
module progmem (
    // Closk & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 10;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin
    mem['h0000] <= 32'h00000093;
    mem['h0001] <= 32'h00000193;
    mem['h0002] <= 32'h00000213;
    mem['h0003] <= 32'h00000293;
    mem['h0004] <= 32'h00000313;
    mem['h0005] <= 32'h00000393;
    mem['h0006] <= 32'h00000413;
    mem['h0007] <= 32'h00000493;
    mem['h0008] <= 32'h00000513;
    mem['h0009] <= 32'h00000593;
    mem['h000A] <= 32'h00000613;
    mem['h000B] <= 32'h00000693;
    mem['h000C] <= 32'h00000713;
    mem['h000D] <= 32'h00000793;
    mem['h000E] <= 32'h00000813;
    mem['h000F] <= 32'h00000893;
    mem['h0010] <= 32'h00000913;
    mem['h0011] <= 32'h00000993;
    mem['h0012] <= 32'h00000A13;
    mem['h0013] <= 32'h00000A93;
    mem['h0014] <= 32'h00000B13;
    mem['h0015] <= 32'h00000B93;
    mem['h0016] <= 32'h00000C13;
    mem['h0017] <= 32'h00000C93;
    mem['h0018] <= 32'h00000D13;
    mem['h0019] <= 32'h00000D93;
    mem['h001A] <= 32'h00000E13;
    mem['h001B] <= 32'h00000E93;
    mem['h001C] <= 32'h00000F13;
    mem['h001D] <= 32'h00000F93;
    mem['h001E] <= 32'h00000513;
    mem['h001F] <= 32'h00000593;
    mem['h0020] <= 32'h00B52023;
    mem['h0021] <= 32'h00450513;
    mem['h0022] <= 32'hFE254CE3;
    mem['h0023] <= 32'h00001517;
    mem['h0024] <= 32'h61050513;
    mem['h0025] <= 32'h00000593;
    mem['h0026] <= 32'h10000613;
    mem['h0027] <= 32'h00C5DC63;
    mem['h0028] <= 32'h00052683;
    mem['h0029] <= 32'h00D5A023;
    mem['h002A] <= 32'h00450513;
    mem['h002B] <= 32'h00458593;
    mem['h002C] <= 32'hFEC5C8E3;
    mem['h002D] <= 32'h10000513;
    mem['h002E] <= 32'h10000593;
    mem['h002F] <= 32'h00B55863;
    mem['h0030] <= 32'h00052023;
    mem['h0031] <= 32'h00450513;
    mem['h0032] <= 32'hFEB54CE3;
    mem['h0033] <= 32'h008000EF;
    mem['h0034] <= 32'h0000006F;
    mem['h0035] <= 32'hFA010113;
    mem['h0036] <= 32'h04112E23;
    mem['h0037] <= 32'h04812C23;
    mem['h0038] <= 32'h06010413;
    mem['h0039] <= 32'h001017B7;
    mem['h003A] <= 32'h65C78793;
    mem['h003B] <= 32'h0007A603;
    mem['h003C] <= 32'h0047A683;
    mem['h003D] <= 32'h0087A703;
    mem['h003E] <= 32'hFEC42023;
    mem['h003F] <= 32'hFED42223;
    mem['h0040] <= 32'hFEE42423;
    mem['h0041] <= 32'h00C7D783;
    mem['h0042] <= 32'hFEF41623;
    mem['h0043] <= 32'h020007B7;
    mem['h0044] <= 32'h00478793;
    mem['h0045] <= 32'h06800713;
    mem['h0046] <= 32'h00E7A023;
    mem['h0047] <= 32'h001017B7;
    mem['h0048] <= 32'h52878513;
    mem['h0049] <= 32'h16C000EF;
    mem['h004A] <= 32'h00000013;
    mem['h004B] <= 32'h001017B7;
    mem['h004C] <= 32'h53C78513;
    mem['h004D] <= 32'h664000EF;
    mem['h004E] <= 32'h00050793;
    mem['h004F] <= 32'h00078713;
    mem['h0050] <= 32'h00D00793;
    mem['h0051] <= 32'hFEF714E3;
    mem['h0052] <= 32'h001017B7;
    mem['h0053] <= 32'h55878513;
    mem['h0054] <= 32'h140000EF;
    mem['h0055] <= 32'h001017B7;
    mem['h0056] <= 32'h55C78513;
    mem['h0057] <= 32'h134000EF;
    mem['h0058] <= 32'h001017B7;
    mem['h0059] <= 32'h58478513;
    mem['h005A] <= 32'h128000EF;
    mem['h005B] <= 32'h001017B7;
    mem['h005C] <= 32'h5AC78513;
    mem['h005D] <= 32'h11C000EF;
    mem['h005E] <= 32'h001017B7;
    mem['h005F] <= 32'h5D078513;
    mem['h0060] <= 32'h110000EF;
    mem['h0061] <= 32'h001017B7;
    mem['h0062] <= 32'h5F878513;
    mem['h0063] <= 32'h104000EF;
    mem['h0064] <= 32'h001017B7;
    mem['h0065] <= 32'h55878513;
    mem['h0066] <= 32'h0F8000EF;
    mem['h0067] <= 32'h001017B7;
    mem['h0068] <= 32'h62078513;
    mem['h0069] <= 32'h0EC000EF;
    mem['h006A] <= 32'hFA040713;
    mem['h006B] <= 32'hFE040793;
    mem['h006C] <= 32'h00070613;
    mem['h006D] <= 32'h00D00593;
    mem['h006E] <= 32'h00078513;
    mem['h006F] <= 32'h284010EF;
    mem['h0070] <= 32'h001017B7;
    mem['h0071] <= 32'h63878513;
    mem['h0072] <= 32'h0C8000EF;
    mem['h0073] <= 32'h001017B7;
    mem['h0074] <= 32'h55878513;
    mem['h0075] <= 32'h0BC000EF;
    mem['h0076] <= 32'h001017B7;
    mem['h0077] <= 32'h64878513;
    mem['h0078] <= 32'h0B0000EF;
    mem['h0079] <= 32'hFE040793;
    mem['h007A] <= 32'h00078513;
    mem['h007B] <= 32'h0A4000EF;
    mem['h007C] <= 32'h001017B7;
    mem['h007D] <= 32'h55878513;
    mem['h007E] <= 32'h098000EF;
    mem['h007F] <= 32'h001017B7;
    mem['h0080] <= 32'h55878513;
    mem['h0081] <= 32'h08C000EF;
    mem['h0082] <= 32'h001017B7;
    mem['h0083] <= 32'h65078513;
    mem['h0084] <= 32'h080000EF;
    mem['h0085] <= 32'hFA040793;
    mem['h0086] <= 32'h00078513;
    mem['h0087] <= 32'h074000EF;
    mem['h0088] <= 32'h001017B7;
    mem['h0089] <= 32'h55878513;
    mem['h008A] <= 32'h068000EF;
    mem['h008B] <= 32'h00000013;
    mem['h008C] <= 32'h05C12083;
    mem['h008D] <= 32'h05812403;
    mem['h008E] <= 32'h06010113;
    mem['h008F] <= 32'h00008067;
    mem['h0090] <= 32'hFE010113;
    mem['h0091] <= 32'h00112E23;
    mem['h0092] <= 32'h00812C23;
    mem['h0093] <= 32'h02010413;
    mem['h0094] <= 32'h00050793;
    mem['h0095] <= 32'hFEF407A3;
    mem['h0096] <= 32'hFEF44703;
    mem['h0097] <= 32'h00A00793;
    mem['h0098] <= 32'h00F71663;
    mem['h0099] <= 32'h00D00513;
    mem['h009A] <= 32'hFD9FF0EF;
    mem['h009B] <= 32'h020007B7;
    mem['h009C] <= 32'h00878793;
    mem['h009D] <= 32'hFEF44703;
    mem['h009E] <= 32'h00E7A023;
    mem['h009F] <= 32'h00000013;
    mem['h00A0] <= 32'h01C12083;
    mem['h00A1] <= 32'h01812403;
    mem['h00A2] <= 32'h02010113;
    mem['h00A3] <= 32'h00008067;
    mem['h00A4] <= 32'hFE010113;
    mem['h00A5] <= 32'h00112E23;
    mem['h00A6] <= 32'h00812C23;
    mem['h00A7] <= 32'h02010413;
    mem['h00A8] <= 32'hFEA42623;
    mem['h00A9] <= 32'h01C0006F;
    mem['h00AA] <= 32'hFEC42783;
    mem['h00AB] <= 32'h00178713;
    mem['h00AC] <= 32'hFEE42623;
    mem['h00AD] <= 32'h0007C783;
    mem['h00AE] <= 32'h00078513;
    mem['h00AF] <= 32'hF85FF0EF;
    mem['h00B0] <= 32'hFEC42783;
    mem['h00B1] <= 32'h0007C783;
    mem['h00B2] <= 32'hFE0790E3;
    mem['h00B3] <= 32'h00000013;
    mem['h00B4] <= 32'h00000013;
    mem['h00B5] <= 32'h01C12083;
    mem['h00B6] <= 32'h01812403;
    mem['h00B7] <= 32'h02010113;
    mem['h00B8] <= 32'h00008067;
    mem['h00B9] <= 32'hFD010113;
    mem['h00BA] <= 32'h02112623;
    mem['h00BB] <= 32'h02812423;
    mem['h00BC] <= 32'h03010413;
    mem['h00BD] <= 32'hFCA42E23;
    mem['h00BE] <= 32'hFCB42C23;
    mem['h00BF] <= 32'h00700793;
    mem['h00C0] <= 32'hFEF42623;
    mem['h00C1] <= 32'h06C0006F;
    mem['h00C2] <= 32'hFEC42783;
    mem['h00C3] <= 32'h00279793;
    mem['h00C4] <= 32'hFDC42703;
    mem['h00C5] <= 32'h00F757B3;
    mem['h00C6] <= 32'h00F7F793;
    mem['h00C7] <= 32'h00101737;
    mem['h00C8] <= 32'h66C70713;
    mem['h00C9] <= 32'h00F707B3;
    mem['h00CA] <= 32'h0007C783;
    mem['h00CB] <= 32'hFEF405A3;
    mem['h00CC] <= 32'hFEB44703;
    mem['h00CD] <= 32'h03000793;
    mem['h00CE] <= 32'h00F71863;
    mem['h00CF] <= 32'hFEC42703;
    mem['h00D0] <= 32'hFD842783;
    mem['h00D1] <= 32'h00F75E63;
    mem['h00D2] <= 32'hFEB44783;
    mem['h00D3] <= 32'h00078513;
    mem['h00D4] <= 32'hEF1FF0EF;
    mem['h00D5] <= 32'hFEC42783;
    mem['h00D6] <= 32'hFCF42C23;
    mem['h00D7] <= 32'h0080006F;
    mem['h00D8] <= 32'h00000013;
    mem['h00D9] <= 32'hFEC42783;
    mem['h00DA] <= 32'hFFF78793;
    mem['h00DB] <= 32'hFEF42623;
    mem['h00DC] <= 32'hFEC42783;
    mem['h00DD] <= 32'hF807DAE3;
    mem['h00DE] <= 32'h00000013;
    mem['h00DF] <= 32'h00000013;
    mem['h00E0] <= 32'h02C12083;
    mem['h00E1] <= 32'h02812403;
    mem['h00E2] <= 32'h03010113;
    mem['h00E3] <= 32'h00008067;
    mem['h00E4] <= 32'hFE010113;
    mem['h00E5] <= 32'h00112E23;
    mem['h00E6] <= 32'h00812C23;
    mem['h00E7] <= 32'h02010413;
    mem['h00E8] <= 32'hFEA42623;
    mem['h00E9] <= 32'hFEC42703;
    mem['h00EA] <= 32'h3E700793;
    mem['h00EB] <= 32'h00E7FA63;
    mem['h00EC] <= 32'h001017B7;
    mem['h00ED] <= 32'h68078513;
    mem['h00EE] <= 32'hED9FF0EF;
    mem['h00EF] <= 32'h3CC0006F;
    mem['h00F0] <= 32'hFEC42703;
    mem['h00F1] <= 32'h38300793;
    mem['h00F2] <= 32'h00E7FE63;
    mem['h00F3] <= 32'h03900513;
    mem['h00F4] <= 32'hE71FF0EF;
    mem['h00F5] <= 32'hFEC42783;
    mem['h00F6] <= 32'hC7C78793;
    mem['h00F7] <= 32'hFEF42623;
    mem['h00F8] <= 32'h1200006F;
    mem['h00F9] <= 32'hFEC42703;
    mem['h00FA] <= 32'h31F00793;
    mem['h00FB] <= 32'h00E7FE63;
    mem['h00FC] <= 32'h03800513;
    mem['h00FD] <= 32'hE4DFF0EF;
    mem['h00FE] <= 32'hFEC42783;
    mem['h00FF] <= 32'hCE078793;
    mem['h0100] <= 32'hFEF42623;
    mem['h0101] <= 32'h0FC0006F;
    mem['h0102] <= 32'hFEC42703;
    mem['h0103] <= 32'h2BB00793;
    mem['h0104] <= 32'h00E7FE63;
    mem['h0105] <= 32'h03700513;
    mem['h0106] <= 32'hE29FF0EF;
    mem['h0107] <= 32'hFEC42783;
    mem['h0108] <= 32'hD4478793;
    mem['h0109] <= 32'hFEF42623;
    mem['h010A] <= 32'h0D80006F;
    mem['h010B] <= 32'hFEC42703;
    mem['h010C] <= 32'h25700793;
    mem['h010D] <= 32'h00E7FE63;
    mem['h010E] <= 32'h03600513;
    mem['h010F] <= 32'hE05FF0EF;
    mem['h0110] <= 32'hFEC42783;
    mem['h0111] <= 32'hDA878793;
    mem['h0112] <= 32'hFEF42623;
    mem['h0113] <= 32'h0B40006F;
    mem['h0114] <= 32'hFEC42703;
    mem['h0115] <= 32'h1F300793;
    mem['h0116] <= 32'h00E7FE63;
    mem['h0117] <= 32'h03500513;
    mem['h0118] <= 32'hDE1FF0EF;
    mem['h0119] <= 32'hFEC42783;
    mem['h011A] <= 32'hE0C78793;
    mem['h011B] <= 32'hFEF42623;
    mem['h011C] <= 32'h0900006F;
    mem['h011D] <= 32'hFEC42703;
    mem['h011E] <= 32'h18F00793;
    mem['h011F] <= 32'h00E7FE63;
    mem['h0120] <= 32'h03400513;
    mem['h0121] <= 32'hDBDFF0EF;
    mem['h0122] <= 32'hFEC42783;
    mem['h0123] <= 32'hE7078793;
    mem['h0124] <= 32'hFEF42623;
    mem['h0125] <= 32'h06C0006F;
    mem['h0126] <= 32'hFEC42703;
    mem['h0127] <= 32'h12B00793;
    mem['h0128] <= 32'h00E7FE63;
    mem['h0129] <= 32'h03300513;
    mem['h012A] <= 32'hD99FF0EF;
    mem['h012B] <= 32'hFEC42783;
    mem['h012C] <= 32'hED478793;
    mem['h012D] <= 32'hFEF42623;
    mem['h012E] <= 32'h0480006F;
    mem['h012F] <= 32'hFEC42703;
    mem['h0130] <= 32'h0C700793;
    mem['h0131] <= 32'h00E7FE63;
    mem['h0132] <= 32'h03200513;
    mem['h0133] <= 32'hD75FF0EF;
    mem['h0134] <= 32'hFEC42783;
    mem['h0135] <= 32'hF3878793;
    mem['h0136] <= 32'hFEF42623;
    mem['h0137] <= 32'h0240006F;
    mem['h0138] <= 32'hFEC42703;
    mem['h0139] <= 32'h06300793;
    mem['h013A] <= 32'h00E7FC63;
    mem['h013B] <= 32'h03100513;
    mem['h013C] <= 32'hD51FF0EF;
    mem['h013D] <= 32'hFEC42783;
    mem['h013E] <= 32'hF9C78793;
    mem['h013F] <= 32'hFEF42623;
    mem['h0140] <= 32'hFEC42703;
    mem['h0141] <= 32'h05900793;
    mem['h0142] <= 32'h00E7FE63;
    mem['h0143] <= 32'h03900513;
    mem['h0144] <= 32'hD31FF0EF;
    mem['h0145] <= 32'hFEC42783;
    mem['h0146] <= 32'hFA678793;
    mem['h0147] <= 32'hFEF42623;
    mem['h0148] <= 32'h1200006F;
    mem['h0149] <= 32'hFEC42703;
    mem['h014A] <= 32'h04F00793;
    mem['h014B] <= 32'h00E7FE63;
    mem['h014C] <= 32'h03800513;
    mem['h014D] <= 32'hD0DFF0EF;
    mem['h014E] <= 32'hFEC42783;
    mem['h014F] <= 32'hFB078793;
    mem['h0150] <= 32'hFEF42623;
    mem['h0151] <= 32'h0FC0006F;
    mem['h0152] <= 32'hFEC42703;
    mem['h0153] <= 32'h04500793;
    mem['h0154] <= 32'h00E7FE63;
    mem['h0155] <= 32'h03700513;
    mem['h0156] <= 32'hCE9FF0EF;
    mem['h0157] <= 32'hFEC42783;
    mem['h0158] <= 32'hFBA78793;
    mem['h0159] <= 32'hFEF42623;
    mem['h015A] <= 32'h0D80006F;
    mem['h015B] <= 32'hFEC42703;
    mem['h015C] <= 32'h03B00793;
    mem['h015D] <= 32'h00E7FE63;
    mem['h015E] <= 32'h03600513;
    mem['h015F] <= 32'hCC5FF0EF;
    mem['h0160] <= 32'hFEC42783;
    mem['h0161] <= 32'hFC478793;
    mem['h0162] <= 32'hFEF42623;
    mem['h0163] <= 32'h0B40006F;
    mem['h0164] <= 32'hFEC42703;
    mem['h0165] <= 32'h03100793;
    mem['h0166] <= 32'h00E7FE63;
    mem['h0167] <= 32'h03500513;
    mem['h0168] <= 32'hCA1FF0EF;
    mem['h0169] <= 32'hFEC42783;
    mem['h016A] <= 32'hFCE78793;
    mem['h016B] <= 32'hFEF42623;
    mem['h016C] <= 32'h0900006F;
    mem['h016D] <= 32'hFEC42703;
    mem['h016E] <= 32'h02700793;
    mem['h016F] <= 32'h00E7FE63;
    mem['h0170] <= 32'h03400513;
    mem['h0171] <= 32'hC7DFF0EF;
    mem['h0172] <= 32'hFEC42783;
    mem['h0173] <= 32'hFD878793;
    mem['h0174] <= 32'hFEF42623;
    mem['h0175] <= 32'h06C0006F;
    mem['h0176] <= 32'hFEC42703;
    mem['h0177] <= 32'h01D00793;
    mem['h0178] <= 32'h00E7FE63;
    mem['h0179] <= 32'h03300513;
    mem['h017A] <= 32'hC59FF0EF;
    mem['h017B] <= 32'hFEC42783;
    mem['h017C] <= 32'hFE278793;
    mem['h017D] <= 32'hFEF42623;
    mem['h017E] <= 32'h0480006F;
    mem['h017F] <= 32'hFEC42703;
    mem['h0180] <= 32'h01300793;
    mem['h0181] <= 32'h00E7FE63;
    mem['h0182] <= 32'h03200513;
    mem['h0183] <= 32'hC35FF0EF;
    mem['h0184] <= 32'hFEC42783;
    mem['h0185] <= 32'hFEC78793;
    mem['h0186] <= 32'hFEF42623;
    mem['h0187] <= 32'h0240006F;
    mem['h0188] <= 32'hFEC42703;
    mem['h0189] <= 32'h00900793;
    mem['h018A] <= 32'h00E7FC63;
    mem['h018B] <= 32'h03100513;
    mem['h018C] <= 32'hC11FF0EF;
    mem['h018D] <= 32'hFEC42783;
    mem['h018E] <= 32'hFF678793;
    mem['h018F] <= 32'hFEF42623;
    mem['h0190] <= 32'hFEC42703;
    mem['h0191] <= 32'h00800793;
    mem['h0192] <= 32'h00E7FE63;
    mem['h0193] <= 32'h03900513;
    mem['h0194] <= 32'hBF1FF0EF;
    mem['h0195] <= 32'hFEC42783;
    mem['h0196] <= 32'hFF778793;
    mem['h0197] <= 32'hFEF42623;
    mem['h0198] <= 32'h1280006F;
    mem['h0199] <= 32'hFEC42703;
    mem['h019A] <= 32'h00700793;
    mem['h019B] <= 32'h00E7FE63;
    mem['h019C] <= 32'h03800513;
    mem['h019D] <= 32'hBCDFF0EF;
    mem['h019E] <= 32'hFEC42783;
    mem['h019F] <= 32'hFF878793;
    mem['h01A0] <= 32'hFEF42623;
    mem['h01A1] <= 32'h1040006F;
    mem['h01A2] <= 32'hFEC42703;
    mem['h01A3] <= 32'h00600793;
    mem['h01A4] <= 32'h00E7FE63;
    mem['h01A5] <= 32'h03700513;
    mem['h01A6] <= 32'hBA9FF0EF;
    mem['h01A7] <= 32'hFEC42783;
    mem['h01A8] <= 32'hFF978793;
    mem['h01A9] <= 32'hFEF42623;
    mem['h01AA] <= 32'h0E00006F;
    mem['h01AB] <= 32'hFEC42703;
    mem['h01AC] <= 32'h00500793;
    mem['h01AD] <= 32'h00E7FE63;
    mem['h01AE] <= 32'h03600513;
    mem['h01AF] <= 32'hB85FF0EF;
    mem['h01B0] <= 32'hFEC42783;
    mem['h01B1] <= 32'hFFA78793;
    mem['h01B2] <= 32'hFEF42623;
    mem['h01B3] <= 32'h0BC0006F;
    mem['h01B4] <= 32'hFEC42703;
    mem['h01B5] <= 32'h00400793;
    mem['h01B6] <= 32'h00E7FE63;
    mem['h01B7] <= 32'h03500513;
    mem['h01B8] <= 32'hB61FF0EF;
    mem['h01B9] <= 32'hFEC42783;
    mem['h01BA] <= 32'hFFB78793;
    mem['h01BB] <= 32'hFEF42623;
    mem['h01BC] <= 32'h0980006F;
    mem['h01BD] <= 32'hFEC42703;
    mem['h01BE] <= 32'h00300793;
    mem['h01BF] <= 32'h00E7FE63;
    mem['h01C0] <= 32'h03400513;
    mem['h01C1] <= 32'hB3DFF0EF;
    mem['h01C2] <= 32'hFEC42783;
    mem['h01C3] <= 32'hFFC78793;
    mem['h01C4] <= 32'hFEF42623;
    mem['h01C5] <= 32'h0740006F;
    mem['h01C6] <= 32'hFEC42703;
    mem['h01C7] <= 32'h00200793;
    mem['h01C8] <= 32'h00E7FE63;
    mem['h01C9] <= 32'h03300513;
    mem['h01CA] <= 32'hB19FF0EF;
    mem['h01CB] <= 32'hFEC42783;
    mem['h01CC] <= 32'hFFD78793;
    mem['h01CD] <= 32'hFEF42623;
    mem['h01CE] <= 32'h0500006F;
    mem['h01CF] <= 32'hFEC42703;
    mem['h01D0] <= 32'h00100793;
    mem['h01D1] <= 32'h00E7FE63;
    mem['h01D2] <= 32'h03200513;
    mem['h01D3] <= 32'hAF5FF0EF;
    mem['h01D4] <= 32'hFEC42783;
    mem['h01D5] <= 32'hFFE78793;
    mem['h01D6] <= 32'hFEF42623;
    mem['h01D7] <= 32'h02C0006F;
    mem['h01D8] <= 32'hFEC42783;
    mem['h01D9] <= 32'h00078E63;
    mem['h01DA] <= 32'h03100513;
    mem['h01DB] <= 32'hAD5FF0EF;
    mem['h01DC] <= 32'hFEC42783;
    mem['h01DD] <= 32'hFFF78793;
    mem['h01DE] <= 32'hFEF42623;
    mem['h01DF] <= 32'h00C0006F;
    mem['h01E0] <= 32'h03000513;
    mem['h01E1] <= 32'hABDFF0EF;
    mem['h01E2] <= 32'h01C12083;
    mem['h01E3] <= 32'h01812403;
    mem['h01E4] <= 32'h02010113;
    mem['h01E5] <= 32'h00008067;
    mem['h01E6] <= 32'hFD010113;
    mem['h01E7] <= 32'h02112623;
    mem['h01E8] <= 32'h02812423;
    mem['h01E9] <= 32'h03010413;
    mem['h01EA] <= 32'hFCA42E23;
    mem['h01EB] <= 32'hFFF00793;
    mem['h01EC] <= 32'hFEF42623;
    mem['h01ED] <= 32'hC00027F3;
    mem['h01EE] <= 32'hFEF42423;
    mem['h01EF] <= 32'hFDC42783;
    mem['h01F0] <= 32'h06078063;
    mem['h01F1] <= 32'hFDC42503;
    mem['h01F2] <= 32'hAC9FF0EF;
    mem['h01F3] <= 32'h0540006F;
    mem['h01F4] <= 32'hC00027F3;
    mem['h01F5] <= 32'hFEF42223;
    mem['h01F6] <= 32'hFE442703;
    mem['h01F7] <= 32'hFE842783;
    mem['h01F8] <= 32'h40F707B3;
    mem['h01F9] <= 32'hFEF42023;
    mem['h01FA] <= 32'hFE042703;
    mem['h01FB] <= 32'h00B727B7;
    mem['h01FC] <= 32'hB0078793;
    mem['h01FD] <= 32'h00E7FE63;
    mem['h01FE] <= 32'hFDC42783;
    mem['h01FF] <= 32'h00078663;
    mem['h0200] <= 32'hFDC42503;
    mem['h0201] <= 32'hA8DFF0EF;
    mem['h0202] <= 32'hFE442783;
    mem['h0203] <= 32'hFEF42423;
    mem['h0204] <= 32'h020007B7;
    mem['h0205] <= 32'h00878793;
    mem['h0206] <= 32'h0007A783;
    mem['h0207] <= 32'hFEF42623;
    mem['h0208] <= 32'hFEC42703;
    mem['h0209] <= 32'hFFF00793;
    mem['h020A] <= 32'hFAF704E3;
    mem['h020B] <= 32'hFEC42783;
    mem['h020C] <= 32'h0FF7F793;
    mem['h020D] <= 32'h00078513;
    mem['h020E] <= 32'h02C12083;
    mem['h020F] <= 32'h02812403;
    mem['h0210] <= 32'h03010113;
    mem['h0211] <= 32'h00008067;
    mem['h0212] <= 32'hFF010113;
    mem['h0213] <= 32'h00112623;
    mem['h0214] <= 32'h00812423;
    mem['h0215] <= 32'h01010413;
    mem['h0216] <= 32'h00000513;
    mem['h0217] <= 32'hF3DFF0EF;
    mem['h0218] <= 32'h00050793;
    mem['h0219] <= 32'h00078513;
    mem['h021A] <= 32'h00C12083;
    mem['h021B] <= 32'h00812403;
    mem['h021C] <= 32'h01010113;
    mem['h021D] <= 32'h00008067;
    mem['h021E] <= 32'hFE010113;
    mem['h021F] <= 32'h00812E23;
    mem['h0220] <= 32'h02010413;
    mem['h0221] <= 32'h00050793;
    mem['h0222] <= 32'hFEB42423;
    mem['h0223] <= 32'hFEF407A3;
    mem['h0224] <= 32'hFEF44783;
    mem['h0225] <= 32'h0047D793;
    mem['h0226] <= 32'h0FF7F793;
    mem['h0227] <= 32'h00F7F793;
    mem['h0228] <= 32'h00101737;
    mem['h0229] <= 32'h68870713;
    mem['h022A] <= 32'h00F707B3;
    mem['h022B] <= 32'h0007C703;
    mem['h022C] <= 32'hFE842783;
    mem['h022D] <= 32'h00E78023;
    mem['h022E] <= 32'hFEF44783;
    mem['h022F] <= 32'h00F7F713;
    mem['h0230] <= 32'hFE842783;
    mem['h0231] <= 32'h00178793;
    mem['h0232] <= 32'h001016B7;
    mem['h0233] <= 32'h68868693;
    mem['h0234] <= 32'h00E68733;
    mem['h0235] <= 32'h00074703;
    mem['h0236] <= 32'h00E78023;
    mem['h0237] <= 32'hFE842783;
    mem['h0238] <= 32'h00278793;
    mem['h0239] <= 32'h00078023;
    mem['h023A] <= 32'h00000013;
    mem['h023B] <= 32'h01C12403;
    mem['h023C] <= 32'h02010113;
    mem['h023D] <= 32'h00008067;
    mem['h023E] <= 32'hF5010113;
    mem['h023F] <= 32'h0A112623;
    mem['h0240] <= 32'h0A812423;
    mem['h0241] <= 32'h0B010413;
    mem['h0242] <= 32'hF4A42E23;
    mem['h0243] <= 32'hF4B42C23;
    mem['h0244] <= 32'hFE042623;
    mem['h0245] <= 32'h0640006F;
    mem['h0246] <= 32'hFEC42783;
    mem['h0247] <= 32'hF5842703;
    mem['h0248] <= 32'h00F707B3;
    mem['h0249] <= 32'h0007C783;
    mem['h024A] <= 32'hF6440713;
    mem['h024B] <= 32'h00070593;
    mem['h024C] <= 32'h00078513;
    mem['h024D] <= 32'hF45FF0EF;
    mem['h024E] <= 32'hFEC42783;
    mem['h024F] <= 32'h00179793;
    mem['h0250] <= 32'hF6444703;
    mem['h0251] <= 32'hFF078793;
    mem['h0252] <= 32'h008787B3;
    mem['h0253] <= 32'hF6E78C23;
    mem['h0254] <= 32'hFEC42783;
    mem['h0255] <= 32'h00179793;
    mem['h0256] <= 32'h00178793;
    mem['h0257] <= 32'hF6544703;
    mem['h0258] <= 32'hFF078793;
    mem['h0259] <= 32'h008787B3;
    mem['h025A] <= 32'hF6E78C23;
    mem['h025B] <= 32'hFEC42783;
    mem['h025C] <= 32'h00178793;
    mem['h025D] <= 32'hFEF42623;
    mem['h025E] <= 32'hFEC42703;
    mem['h025F] <= 32'h03F00793;
    mem['h0260] <= 32'hF8E7DCE3;
    mem['h0261] <= 32'hFE040423;
    mem['h0262] <= 32'h00000013;
    mem['h0263] <= 32'h0AC12083;
    mem['h0264] <= 32'h0A812403;
    mem['h0265] <= 32'h0B010113;
    mem['h0266] <= 32'h00008067;
    mem['h0267] <= 32'hEB010113;
    mem['h0268] <= 32'h14812623;
    mem['h0269] <= 32'h15010413;
    mem['h026A] <= 32'hEAA42E23;
    mem['h026B] <= 32'hEAB42C23;
    mem['h026C] <= 32'hFC042623;
    mem['h026D] <= 32'hFC042423;
    mem['h026E] <= 32'h0980006F;
    mem['h026F] <= 32'hEB842703;
    mem['h0270] <= 32'hFC842783;
    mem['h0271] <= 32'h00F707B3;
    mem['h0272] <= 32'h0007C783;
    mem['h0273] <= 32'h01879713;
    mem['h0274] <= 32'hFC842783;
    mem['h0275] <= 32'h00178793;
    mem['h0276] <= 32'hEB842683;
    mem['h0277] <= 32'h00F687B3;
    mem['h0278] <= 32'h0007C783;
    mem['h0279] <= 32'h01079793;
    mem['h027A] <= 32'h00F76733;
    mem['h027B] <= 32'hFC842783;
    mem['h027C] <= 32'h00278793;
    mem['h027D] <= 32'hEB842683;
    mem['h027E] <= 32'h00F687B3;
    mem['h027F] <= 32'h0007C783;
    mem['h0280] <= 32'h00879793;
    mem['h0281] <= 32'h00F767B3;
    mem['h0282] <= 32'hFC842703;
    mem['h0283] <= 32'h00370713;
    mem['h0284] <= 32'hEB842683;
    mem['h0285] <= 32'h00E68733;
    mem['h0286] <= 32'h00074703;
    mem['h0287] <= 32'h00E7E7B3;
    mem['h0288] <= 32'h00078713;
    mem['h0289] <= 32'hFCC42783;
    mem['h028A] <= 32'h00279793;
    mem['h028B] <= 32'hFF078793;
    mem['h028C] <= 32'h008787B3;
    mem['h028D] <= 32'hECE7A823;
    mem['h028E] <= 32'hFCC42783;
    mem['h028F] <= 32'h00178793;
    mem['h0290] <= 32'hFCF42623;
    mem['h0291] <= 32'hFC842783;
    mem['h0292] <= 32'h00478793;
    mem['h0293] <= 32'hFCF42423;
    mem['h0294] <= 32'hFCC42703;
    mem['h0295] <= 32'h00F00793;
    mem['h0296] <= 32'hF6E7F2E3;
    mem['h0297] <= 32'h1380006F;
    mem['h0298] <= 32'hFCC42783;
    mem['h0299] <= 32'hFFE78793;
    mem['h029A] <= 32'h00279793;
    mem['h029B] <= 32'hFF078793;
    mem['h029C] <= 32'h008787B3;
    mem['h029D] <= 32'hED07A783;
    mem['h029E] <= 32'h00F79693;
    mem['h029F] <= 32'h0117D713;
    mem['h02A0] <= 32'h00D76733;
    mem['h02A1] <= 32'hFCC42783;
    mem['h02A2] <= 32'hFFE78793;
    mem['h02A3] <= 32'h00279793;
    mem['h02A4] <= 32'hFF078793;
    mem['h02A5] <= 32'h008787B3;
    mem['h02A6] <= 32'hED07A783;
    mem['h02A7] <= 32'h00D79693;
    mem['h02A8] <= 32'h0137D793;
    mem['h02A9] <= 32'h00D7E7B3;
    mem['h02AA] <= 32'h00F74733;
    mem['h02AB] <= 32'hFCC42783;
    mem['h02AC] <= 32'hFFE78793;
    mem['h02AD] <= 32'h00279793;
    mem['h02AE] <= 32'hFF078793;
    mem['h02AF] <= 32'h008787B3;
    mem['h02B0] <= 32'hED07A783;
    mem['h02B1] <= 32'h00A7D793;
    mem['h02B2] <= 32'h00F74733;
    mem['h02B3] <= 32'hFCC42783;
    mem['h02B4] <= 32'hFF978793;
    mem['h02B5] <= 32'h00279793;
    mem['h02B6] <= 32'hFF078793;
    mem['h02B7] <= 32'h008787B3;
    mem['h02B8] <= 32'hED07A783;
    mem['h02B9] <= 32'h00F706B3;
    mem['h02BA] <= 32'hFCC42783;
    mem['h02BB] <= 32'hFF178793;
    mem['h02BC] <= 32'h00279793;
    mem['h02BD] <= 32'hFF078793;
    mem['h02BE] <= 32'h008787B3;
    mem['h02BF] <= 32'hED07A783;
    mem['h02C0] <= 32'h0077D613;
    mem['h02C1] <= 32'h01979713;
    mem['h02C2] <= 32'h00C76733;
    mem['h02C3] <= 32'hFCC42783;
    mem['h02C4] <= 32'hFF178793;
    mem['h02C5] <= 32'h00279793;
    mem['h02C6] <= 32'hFF078793;
    mem['h02C7] <= 32'h008787B3;
    mem['h02C8] <= 32'hED07A783;
    mem['h02C9] <= 32'h00E79613;
    mem['h02CA] <= 32'h0127D793;
    mem['h02CB] <= 32'h00C7E7B3;
    mem['h02CC] <= 32'h00F74733;
    mem['h02CD] <= 32'hFCC42783;
    mem['h02CE] <= 32'hFF178793;
    mem['h02CF] <= 32'h00279793;
    mem['h02D0] <= 32'hFF078793;
    mem['h02D1] <= 32'h008787B3;
    mem['h02D2] <= 32'hED07A783;
    mem['h02D3] <= 32'h0037D793;
    mem['h02D4] <= 32'h00F747B3;
    mem['h02D5] <= 32'h00F68733;
    mem['h02D6] <= 32'hFCC42783;
    mem['h02D7] <= 32'hFF078793;
    mem['h02D8] <= 32'h00279793;
    mem['h02D9] <= 32'hFF078793;
    mem['h02DA] <= 32'h008787B3;
    mem['h02DB] <= 32'hED07A783;
    mem['h02DC] <= 32'h00F70733;
    mem['h02DD] <= 32'hFCC42783;
    mem['h02DE] <= 32'h00279793;
    mem['h02DF] <= 32'hFF078793;
    mem['h02E0] <= 32'h008787B3;
    mem['h02E1] <= 32'hECE7A823;
    mem['h02E2] <= 32'hFCC42783;
    mem['h02E3] <= 32'h00178793;
    mem['h02E4] <= 32'hFCF42623;
    mem['h02E5] <= 32'hFCC42703;
    mem['h02E6] <= 32'h03F00793;
    mem['h02E7] <= 32'hECE7F2E3;
    mem['h02E8] <= 32'hEBC42783;
    mem['h02E9] <= 32'h0507A783;
    mem['h02EA] <= 32'hFEF42623;
    mem['h02EB] <= 32'hEBC42783;
    mem['h02EC] <= 32'h0547A783;
    mem['h02ED] <= 32'hFEF42423;
    mem['h02EE] <= 32'hEBC42783;
    mem['h02EF] <= 32'h0587A783;
    mem['h02F0] <= 32'hFEF42223;
    mem['h02F1] <= 32'hEBC42783;
    mem['h02F2] <= 32'h05C7A783;
    mem['h02F3] <= 32'hFEF42023;
    mem['h02F4] <= 32'hEBC42783;
    mem['h02F5] <= 32'h0607A783;
    mem['h02F6] <= 32'hFCF42E23;
    mem['h02F7] <= 32'hEBC42783;
    mem['h02F8] <= 32'h0647A783;
    mem['h02F9] <= 32'hFCF42C23;
    mem['h02FA] <= 32'hEBC42783;
    mem['h02FB] <= 32'h0687A783;
    mem['h02FC] <= 32'hFCF42A23;
    mem['h02FD] <= 32'hEBC42783;
    mem['h02FE] <= 32'h06C7A783;
    mem['h02FF] <= 32'hFCF42823;
    mem['h0300] <= 32'hFC042623;
    mem['h0301] <= 32'h15C0006F;
    mem['h0302] <= 32'hFDC42783;
    mem['h0303] <= 32'h0067D693;
    mem['h0304] <= 32'h01A79713;
    mem['h0305] <= 32'h00D76733;
    mem['h0306] <= 32'hFDC42783;
    mem['h0307] <= 32'h00B7D693;
    mem['h0308] <= 32'h01579793;
    mem['h0309] <= 32'h00D7E7B3;
    mem['h030A] <= 32'h00F74733;
    mem['h030B] <= 32'hFDC42783;
    mem['h030C] <= 32'h00779693;
    mem['h030D] <= 32'h0197D793;
    mem['h030E] <= 32'h00D7E7B3;
    mem['h030F] <= 32'h00F74733;
    mem['h0310] <= 32'hFD042783;
    mem['h0311] <= 32'h00F70733;
    mem['h0312] <= 32'hFDC42683;
    mem['h0313] <= 32'hFD842783;
    mem['h0314] <= 32'h00F6F6B3;
    mem['h0315] <= 32'hFDC42783;
    mem['h0316] <= 32'hFFF7C613;
    mem['h0317] <= 32'hFD442783;
    mem['h0318] <= 32'h00F677B3;
    mem['h0319] <= 32'h00F6C7B3;
    mem['h031A] <= 32'h00F70733;
    mem['h031B] <= 32'h00000693;
    mem['h031C] <= 32'hFCC42783;
    mem['h031D] <= 32'h00279793;
    mem['h031E] <= 32'h00F687B3;
    mem['h031F] <= 32'h0007A783;
    mem['h0320] <= 32'h00F70733;
    mem['h0321] <= 32'hFCC42783;
    mem['h0322] <= 32'h00279793;
    mem['h0323] <= 32'hFF078793;
    mem['h0324] <= 32'h008787B3;
    mem['h0325] <= 32'hED07A783;
    mem['h0326] <= 32'h00F707B3;
    mem['h0327] <= 32'hFCF42223;
    mem['h0328] <= 32'hFEC42783;
    mem['h0329] <= 32'h0027D693;
    mem['h032A] <= 32'h01E79713;
    mem['h032B] <= 32'h00D76733;
    mem['h032C] <= 32'hFEC42783;
    mem['h032D] <= 32'h00D7D693;
    mem['h032E] <= 32'h01379793;
    mem['h032F] <= 32'h00D7E7B3;
    mem['h0330] <= 32'h00F74733;
    mem['h0331] <= 32'hFEC42783;
    mem['h0332] <= 32'h00A79693;
    mem['h0333] <= 32'h0167D793;
    mem['h0334] <= 32'h00D7E7B3;
    mem['h0335] <= 32'h00F74733;
    mem['h0336] <= 32'hFE842683;
    mem['h0337] <= 32'hFE442783;
    mem['h0338] <= 32'h00F6C6B3;
    mem['h0339] <= 32'hFEC42783;
    mem['h033A] <= 32'h00F6F6B3;
    mem['h033B] <= 32'hFE842603;
    mem['h033C] <= 32'hFE442783;
    mem['h033D] <= 32'h00F677B3;
    mem['h033E] <= 32'h00F6C7B3;
    mem['h033F] <= 32'h00F707B3;
    mem['h0340] <= 32'hFCF42023;
    mem['h0341] <= 32'hFD442783;
    mem['h0342] <= 32'hFCF42823;
    mem['h0343] <= 32'hFD842783;
    mem['h0344] <= 32'hFCF42A23;
    mem['h0345] <= 32'hFDC42783;
    mem['h0346] <= 32'hFCF42C23;
    mem['h0347] <= 32'hFE042703;
    mem['h0348] <= 32'hFC442783;
    mem['h0349] <= 32'h00F707B3;
    mem['h034A] <= 32'hFCF42E23;
    mem['h034B] <= 32'hFE442783;
    mem['h034C] <= 32'hFEF42023;
    mem['h034D] <= 32'hFE842783;
    mem['h034E] <= 32'hFEF42223;
    mem['h034F] <= 32'hFEC42783;
    mem['h0350] <= 32'hFEF42423;
    mem['h0351] <= 32'hFC442703;
    mem['h0352] <= 32'hFC042783;
    mem['h0353] <= 32'h00F707B3;
    mem['h0354] <= 32'hFEF42623;
    mem['h0355] <= 32'hFCC42783;
    mem['h0356] <= 32'h00178793;
    mem['h0357] <= 32'hFCF42623;
    mem['h0358] <= 32'hFCC42703;
    mem['h0359] <= 32'h03F00793;
    mem['h035A] <= 32'hEAE7F0E3;
    mem['h035B] <= 32'hEBC42783;
    mem['h035C] <= 32'h0507A703;
    mem['h035D] <= 32'hFEC42783;
    mem['h035E] <= 32'h00F70733;
    mem['h035F] <= 32'hEBC42783;
    mem['h0360] <= 32'h04E7A823;
    mem['h0361] <= 32'hEBC42783;
    mem['h0362] <= 32'h0547A703;
    mem['h0363] <= 32'hFE842783;
    mem['h0364] <= 32'h00F70733;
    mem['h0365] <= 32'hEBC42783;
    mem['h0366] <= 32'h04E7AA23;
    mem['h0367] <= 32'hEBC42783;
    mem['h0368] <= 32'h0587A703;
    mem['h0369] <= 32'hFE442783;
    mem['h036A] <= 32'h00F70733;
    mem['h036B] <= 32'hEBC42783;
    mem['h036C] <= 32'h04E7AC23;
    mem['h036D] <= 32'hEBC42783;
    mem['h036E] <= 32'h05C7A703;
    mem['h036F] <= 32'hFE042783;
    mem['h0370] <= 32'h00F70733;
    mem['h0371] <= 32'hEBC42783;
    mem['h0372] <= 32'h04E7AE23;
    mem['h0373] <= 32'hEBC42783;
    mem['h0374] <= 32'h0607A703;
    mem['h0375] <= 32'hFDC42783;
    mem['h0376] <= 32'h00F70733;
    mem['h0377] <= 32'hEBC42783;
    mem['h0378] <= 32'h06E7A023;
    mem['h0379] <= 32'hEBC42783;
    mem['h037A] <= 32'h0647A703;
    mem['h037B] <= 32'hFD842783;
    mem['h037C] <= 32'h00F70733;
    mem['h037D] <= 32'hEBC42783;
    mem['h037E] <= 32'h06E7A223;
    mem['h037F] <= 32'hEBC42783;
    mem['h0380] <= 32'h0687A703;
    mem['h0381] <= 32'hFD442783;
    mem['h0382] <= 32'h00F70733;
    mem['h0383] <= 32'hEBC42783;
    mem['h0384] <= 32'h06E7A423;
    mem['h0385] <= 32'hEBC42783;
    mem['h0386] <= 32'h06C7A703;
    mem['h0387] <= 32'hFD042783;
    mem['h0388] <= 32'h00F70733;
    mem['h0389] <= 32'hEBC42783;
    mem['h038A] <= 32'h06E7A623;
    mem['h038B] <= 32'h00000013;
    mem['h038C] <= 32'h14C12403;
    mem['h038D] <= 32'h15010113;
    mem['h038E] <= 32'h00008067;
    mem['h038F] <= 32'hFE010113;
    mem['h0390] <= 32'h00812E23;
    mem['h0391] <= 32'h02010413;
    mem['h0392] <= 32'hFEA42623;
    mem['h0393] <= 32'hFEC42783;
    mem['h0394] <= 32'h0407A023;
    mem['h0395] <= 32'hFEC42783;
    mem['h0396] <= 32'h0407A223;
    mem['h0397] <= 32'hFEC42783;
    mem['h0398] <= 32'h0407A423;
    mem['h0399] <= 32'hFEC42783;
    mem['h039A] <= 32'h0407A623;
    mem['h039B] <= 32'hFEC42783;
    mem['h039C] <= 32'h6A09E737;
    mem['h039D] <= 32'h66770713;
    mem['h039E] <= 32'h04E7A823;
    mem['h039F] <= 32'hFEC42783;
    mem['h03A0] <= 32'hBB67B737;
    mem['h03A1] <= 32'hE8570713;
    mem['h03A2] <= 32'h04E7AA23;
    mem['h03A3] <= 32'hFEC42783;
    mem['h03A4] <= 32'h3C6EF737;
    mem['h03A5] <= 32'h37270713;
    mem['h03A6] <= 32'h04E7AC23;
    mem['h03A7] <= 32'hFEC42783;
    mem['h03A8] <= 32'hA54FF737;
    mem['h03A9] <= 32'h53A70713;
    mem['h03AA] <= 32'h04E7AE23;
    mem['h03AB] <= 32'hFEC42783;
    mem['h03AC] <= 32'h510E5737;
    mem['h03AD] <= 32'h27F70713;
    mem['h03AE] <= 32'h06E7A023;
    mem['h03AF] <= 32'hFEC42783;
    mem['h03B0] <= 32'h9B057737;
    mem['h03B1] <= 32'h88C70713;
    mem['h03B2] <= 32'h06E7A223;
    mem['h03B3] <= 32'hFEC42783;
    mem['h03B4] <= 32'h1F83E737;
    mem['h03B5] <= 32'h9AB70713;
    mem['h03B6] <= 32'h06E7A423;
    mem['h03B7] <= 32'hFEC42783;
    mem['h03B8] <= 32'h5BE0D737;
    mem['h03B9] <= 32'hD1970713;
    mem['h03BA] <= 32'h06E7A623;
    mem['h03BB] <= 32'h00000013;
    mem['h03BC] <= 32'h01C12403;
    mem['h03BD] <= 32'h02010113;
    mem['h03BE] <= 32'h00008067;
    mem['h03BF] <= 32'hFD010113;
    mem['h03C0] <= 32'h02112623;
    mem['h03C1] <= 32'h02812423;
    mem['h03C2] <= 32'h03010413;
    mem['h03C3] <= 32'hFCA42E23;
    mem['h03C4] <= 32'hFCB42C23;
    mem['h03C5] <= 32'hFCC42A23;
    mem['h03C6] <= 32'hFE042623;
    mem['h03C7] <= 32'h0CC0006F;
    mem['h03C8] <= 32'hFEC42783;
    mem['h03C9] <= 32'hFD842703;
    mem['h03CA] <= 32'h00F70733;
    mem['h03CB] <= 32'hFDC42783;
    mem['h03CC] <= 32'h0407A783;
    mem['h03CD] <= 32'h00074703;
    mem['h03CE] <= 32'hFDC42683;
    mem['h03CF] <= 32'h00F687B3;
    mem['h03D0] <= 32'h00E78023;
    mem['h03D1] <= 32'hFDC42783;
    mem['h03D2] <= 32'h0407A783;
    mem['h03D3] <= 32'h00178713;
    mem['h03D4] <= 32'hFDC42783;
    mem['h03D5] <= 32'h04E7A023;
    mem['h03D6] <= 32'hFDC42783;
    mem['h03D7] <= 32'h0407A703;
    mem['h03D8] <= 32'h04000793;
    mem['h03D9] <= 32'h06F71C63;
    mem['h03DA] <= 32'hFDC42783;
    mem['h03DB] <= 32'h0447A783;
    mem['h03DC] <= 32'h00178713;
    mem['h03DD] <= 32'hFDC42783;
    mem['h03DE] <= 32'h04E7A223;
    mem['h03DF] <= 32'hFDC42783;
    mem['h03E0] <= 32'h00078593;
    mem['h03E1] <= 32'hFDC42503;
    mem['h03E2] <= 32'h971FF0EF;
    mem['h03E3] <= 32'hFDC42783;
    mem['h03E4] <= 32'h00078593;
    mem['h03E5] <= 32'hFDC42503;
    mem['h03E6] <= 32'hA05FF0EF;
    mem['h03E7] <= 32'hFDC42783;
    mem['h03E8] <= 32'h0487A703;
    mem['h03E9] <= 32'hDFF00793;
    mem['h03EA] <= 32'h00E7FC63;
    mem['h03EB] <= 32'hFDC42783;
    mem['h03EC] <= 32'h04C7A783;
    mem['h03ED] <= 32'h00178713;
    mem['h03EE] <= 32'hFDC42783;
    mem['h03EF] <= 32'h04E7A623;
    mem['h03F0] <= 32'hFDC42783;
    mem['h03F1] <= 32'h0487A783;
    mem['h03F2] <= 32'h20078713;
    mem['h03F3] <= 32'hFDC42783;
    mem['h03F4] <= 32'h04E7A423;
    mem['h03F5] <= 32'hFDC42783;
    mem['h03F6] <= 32'h0407A023;
    mem['h03F7] <= 32'hFEC42783;
    mem['h03F8] <= 32'h00178793;
    mem['h03F9] <= 32'hFEF42623;
    mem['h03FA] <= 32'hFEC42783;
    mem['h03FB] <= 32'hFD442703;
    mem['h03FC] <= 32'hF2E7E8E3;
    mem['h03FD] <= 32'h00000013;
    mem['h03FE] <= 32'h00000013;
    mem['h03FF] <= 32'h02C12083;
    mem['h0400] <= 32'h02812403;
    mem['h0401] <= 32'h03010113;
    mem['h0402] <= 32'h00008067;
    mem['h0403] <= 32'hFD010113;
    mem['h0404] <= 32'h02112623;
    mem['h0405] <= 32'h02812423;
    mem['h0406] <= 32'h03010413;
    mem['h0407] <= 32'hFCA42E23;
    mem['h0408] <= 32'hFCB42C23;
    mem['h0409] <= 32'hFDC42783;
    mem['h040A] <= 32'h0407A783;
    mem['h040B] <= 32'hFEF42623;
    mem['h040C] <= 32'hFDC42783;
    mem['h040D] <= 32'h0407A703;
    mem['h040E] <= 32'h03700793;
    mem['h040F] <= 32'h04E7E663;
    mem['h0410] <= 32'hFEC42783;
    mem['h0411] <= 32'h00178713;
    mem['h0412] <= 32'hFEE42623;
    mem['h0413] <= 32'hFDC42703;
    mem['h0414] <= 32'h00F707B3;
    mem['h0415] <= 32'hF8000713;
    mem['h0416] <= 32'h00E78023;
    mem['h0417] <= 32'h01C0006F;
    mem['h0418] <= 32'hFEC42783;
    mem['h0419] <= 32'h00178713;
    mem['h041A] <= 32'hFEE42623;
    mem['h041B] <= 32'hFDC42703;
    mem['h041C] <= 32'h00F707B3;
    mem['h041D] <= 32'h00078023;
    mem['h041E] <= 32'hFEC42703;
    mem['h041F] <= 32'h03700793;
    mem['h0420] <= 32'hFEE7D0E3;
    mem['h0421] <= 32'h0AC0006F;
    mem['h0422] <= 32'hFEC42783;
    mem['h0423] <= 32'h00178713;
    mem['h0424] <= 32'hFEE42623;
    mem['h0425] <= 32'hFDC42703;
    mem['h0426] <= 32'h00F707B3;
    mem['h0427] <= 32'hF8000713;
    mem['h0428] <= 32'h00E78023;
    mem['h0429] <= 32'h01C0006F;
    mem['h042A] <= 32'hFEC42783;
    mem['h042B] <= 32'h00178713;
    mem['h042C] <= 32'hFEE42623;
    mem['h042D] <= 32'hFDC42703;
    mem['h042E] <= 32'h00F707B3;
    mem['h042F] <= 32'h00078023;
    mem['h0430] <= 32'hFEC42703;
    mem['h0431] <= 32'h03F00793;
    mem['h0432] <= 32'hFEE7D0E3;
    mem['h0433] <= 32'hFDC42783;
    mem['h0434] <= 32'h0447A783;
    mem['h0435] <= 32'h00178713;
    mem['h0436] <= 32'hFDC42783;
    mem['h0437] <= 32'h04E7A223;
    mem['h0438] <= 32'hFDC42783;
    mem['h0439] <= 32'h00078593;
    mem['h043A] <= 32'hFDC42503;
    mem['h043B] <= 32'h80DFF0EF;
    mem['h043C] <= 32'hFDC42783;
    mem['h043D] <= 32'h00078593;
    mem['h043E] <= 32'hFDC42503;
    mem['h043F] <= 32'h8A1FF0EF;
    mem['h0440] <= 32'hFE042423;
    mem['h0441] <= 32'h0200006F;
    mem['h0442] <= 32'hFDC42703;
    mem['h0443] <= 32'hFE842783;
    mem['h0444] <= 32'h00F707B3;
    mem['h0445] <= 32'h00078023;
    mem['h0446] <= 32'hFE842783;
    mem['h0447] <= 32'h00178793;
    mem['h0448] <= 32'hFEF42423;
    mem['h0449] <= 32'hFE842703;
    mem['h044A] <= 32'h03700793;
    mem['h044B] <= 32'hFCE7DEE3;
    mem['h044C] <= 32'hFDC42783;
    mem['h044D] <= 32'h0487A703;
    mem['h044E] <= 32'hFDC42783;
    mem['h044F] <= 32'h0407A783;
    mem['h0450] <= 32'h00379793;
    mem['h0451] <= 32'hFFF7C793;
    mem['h0452] <= 32'h00E7FC63;
    mem['h0453] <= 32'hFDC42783;
    mem['h0454] <= 32'h04C7A783;
    mem['h0455] <= 32'h00178713;
    mem['h0456] <= 32'hFDC42783;
    mem['h0457] <= 32'h04E7A623;
    mem['h0458] <= 32'hFDC42783;
    mem['h0459] <= 32'h0487A703;
    mem['h045A] <= 32'hFDC42783;
    mem['h045B] <= 32'h0407A783;
    mem['h045C] <= 32'h00379793;
    mem['h045D] <= 32'h00F70733;
    mem['h045E] <= 32'hFDC42783;
    mem['h045F] <= 32'h04E7A423;
    mem['h0460] <= 32'hFDC42783;
    mem['h0461] <= 32'h0487A783;
    mem['h0462] <= 32'h0FF7F713;
    mem['h0463] <= 32'hFDC42783;
    mem['h0464] <= 32'h02E78FA3;
    mem['h0465] <= 32'hFDC42783;
    mem['h0466] <= 32'h0487A783;
    mem['h0467] <= 32'h0087D793;
    mem['h0468] <= 32'h0FF7F713;
    mem['h0469] <= 32'hFDC42783;
    mem['h046A] <= 32'h02E78F23;
    mem['h046B] <= 32'hFDC42783;
    mem['h046C] <= 32'h0487A783;
    mem['h046D] <= 32'h0107D793;
    mem['h046E] <= 32'h0FF7F713;
    mem['h046F] <= 32'hFDC42783;
    mem['h0470] <= 32'h02E78EA3;
    mem['h0471] <= 32'hFDC42783;
    mem['h0472] <= 32'h0487A783;
    mem['h0473] <= 32'h0187D793;
    mem['h0474] <= 32'h0FF7F713;
    mem['h0475] <= 32'hFDC42783;
    mem['h0476] <= 32'h02E78E23;
    mem['h0477] <= 32'hFDC42783;
    mem['h0478] <= 32'h04C7A783;
    mem['h0479] <= 32'h0FF7F713;
    mem['h047A] <= 32'hFDC42783;
    mem['h047B] <= 32'h02E78DA3;
    mem['h047C] <= 32'hFDC42783;
    mem['h047D] <= 32'h04C7A783;
    mem['h047E] <= 32'h0087D793;
    mem['h047F] <= 32'h0FF7F713;
    mem['h0480] <= 32'hFDC42783;
    mem['h0481] <= 32'h02E78D23;
    mem['h0482] <= 32'hFDC42783;
    mem['h0483] <= 32'h04C7A783;
    mem['h0484] <= 32'h0107D793;
    mem['h0485] <= 32'h0FF7F713;
    mem['h0486] <= 32'hFDC42783;
    mem['h0487] <= 32'h02E78CA3;
    mem['h0488] <= 32'hFDC42783;
    mem['h0489] <= 32'h04C7A783;
    mem['h048A] <= 32'h0187D793;
    mem['h048B] <= 32'h0FF7F713;
    mem['h048C] <= 32'hFDC42783;
    mem['h048D] <= 32'h02E78C23;
    mem['h048E] <= 32'hFDC42783;
    mem['h048F] <= 32'h0447A783;
    mem['h0490] <= 32'h00178713;
    mem['h0491] <= 32'hFDC42783;
    mem['h0492] <= 32'h04E7A223;
    mem['h0493] <= 32'hFDC42783;
    mem['h0494] <= 32'h00078593;
    mem['h0495] <= 32'hFDC42503;
    mem['h0496] <= 32'hEA0FF0EF;
    mem['h0497] <= 32'hFDC42783;
    mem['h0498] <= 32'h00078593;
    mem['h0499] <= 32'hFDC42503;
    mem['h049A] <= 32'hF34FF0EF;
    mem['h049B] <= 32'hFE042623;
    mem['h049C] <= 32'h1AC0006F;
    mem['h049D] <= 32'hFDC42783;
    mem['h049E] <= 32'h0507A703;
    mem['h049F] <= 32'h00300693;
    mem['h04A0] <= 32'hFEC42783;
    mem['h04A1] <= 32'h40F687B3;
    mem['h04A2] <= 32'h00379793;
    mem['h04A3] <= 32'h00F756B3;
    mem['h04A4] <= 32'hFEC42783;
    mem['h04A5] <= 32'hFD842703;
    mem['h04A6] <= 32'h00F707B3;
    mem['h04A7] <= 32'h0FF6F713;
    mem['h04A8] <= 32'h00E78023;
    mem['h04A9] <= 32'hFDC42783;
    mem['h04AA] <= 32'h0547A703;
    mem['h04AB] <= 32'h00300693;
    mem['h04AC] <= 32'hFEC42783;
    mem['h04AD] <= 32'h40F687B3;
    mem['h04AE] <= 32'h00379793;
    mem['h04AF] <= 32'h00F756B3;
    mem['h04B0] <= 32'hFEC42783;
    mem['h04B1] <= 32'h00478793;
    mem['h04B2] <= 32'hFD842703;
    mem['h04B3] <= 32'h00F707B3;
    mem['h04B4] <= 32'h0FF6F713;
    mem['h04B5] <= 32'h00E78023;
    mem['h04B6] <= 32'hFDC42783;
    mem['h04B7] <= 32'h0587A703;
    mem['h04B8] <= 32'h00300693;
    mem['h04B9] <= 32'hFEC42783;
    mem['h04BA] <= 32'h40F687B3;
    mem['h04BB] <= 32'h00379793;
    mem['h04BC] <= 32'h00F756B3;
    mem['h04BD] <= 32'hFEC42783;
    mem['h04BE] <= 32'h00878793;
    mem['h04BF] <= 32'hFD842703;
    mem['h04C0] <= 32'h00F707B3;
    mem['h04C1] <= 32'h0FF6F713;
    mem['h04C2] <= 32'h00E78023;
    mem['h04C3] <= 32'hFDC42783;
    mem['h04C4] <= 32'h05C7A703;
    mem['h04C5] <= 32'h00300693;
    mem['h04C6] <= 32'hFEC42783;
    mem['h04C7] <= 32'h40F687B3;
    mem['h04C8] <= 32'h00379793;
    mem['h04C9] <= 32'h00F756B3;
    mem['h04CA] <= 32'hFEC42783;
    mem['h04CB] <= 32'h00C78793;
    mem['h04CC] <= 32'hFD842703;
    mem['h04CD] <= 32'h00F707B3;
    mem['h04CE] <= 32'h0FF6F713;
    mem['h04CF] <= 32'h00E78023;
    mem['h04D0] <= 32'hFDC42783;
    mem['h04D1] <= 32'h0607A703;
    mem['h04D2] <= 32'h00300693;
    mem['h04D3] <= 32'hFEC42783;
    mem['h04D4] <= 32'h40F687B3;
    mem['h04D5] <= 32'h00379793;
    mem['h04D6] <= 32'h00F756B3;
    mem['h04D7] <= 32'hFEC42783;
    mem['h04D8] <= 32'h01078793;
    mem['h04D9] <= 32'hFD842703;
    mem['h04DA] <= 32'h00F707B3;
    mem['h04DB] <= 32'h0FF6F713;
    mem['h04DC] <= 32'h00E78023;
    mem['h04DD] <= 32'hFDC42783;
    mem['h04DE] <= 32'h0647A703;
    mem['h04DF] <= 32'h00300693;
    mem['h04E0] <= 32'hFEC42783;
    mem['h04E1] <= 32'h40F687B3;
    mem['h04E2] <= 32'h00379793;
    mem['h04E3] <= 32'h00F756B3;
    mem['h04E4] <= 32'hFEC42783;
    mem['h04E5] <= 32'h01478793;
    mem['h04E6] <= 32'hFD842703;
    mem['h04E7] <= 32'h00F707B3;
    mem['h04E8] <= 32'h0FF6F713;
    mem['h04E9] <= 32'h00E78023;
    mem['h04EA] <= 32'hFDC42783;
    mem['h04EB] <= 32'h0687A703;
    mem['h04EC] <= 32'h00300693;
    mem['h04ED] <= 32'hFEC42783;
    mem['h04EE] <= 32'h40F687B3;
    mem['h04EF] <= 32'h00379793;
    mem['h04F0] <= 32'h00F756B3;
    mem['h04F1] <= 32'hFEC42783;
    mem['h04F2] <= 32'h01878793;
    mem['h04F3] <= 32'hFD842703;
    mem['h04F4] <= 32'h00F707B3;
    mem['h04F5] <= 32'h0FF6F713;
    mem['h04F6] <= 32'h00E78023;
    mem['h04F7] <= 32'hFDC42783;
    mem['h04F8] <= 32'h06C7A703;
    mem['h04F9] <= 32'h00300693;
    mem['h04FA] <= 32'hFEC42783;
    mem['h04FB] <= 32'h40F687B3;
    mem['h04FC] <= 32'h00379793;
    mem['h04FD] <= 32'h00F756B3;
    mem['h04FE] <= 32'hFEC42783;
    mem['h04FF] <= 32'h01C78793;
    mem['h0500] <= 32'hFD842703;
    mem['h0501] <= 32'h00F707B3;
    mem['h0502] <= 32'h0FF6F713;
    mem['h0503] <= 32'h00E78023;
    mem['h0504] <= 32'hFEC42783;
    mem['h0505] <= 32'h00178793;
    mem['h0506] <= 32'hFEF42623;
    mem['h0507] <= 32'hFEC42703;
    mem['h0508] <= 32'h00300793;
    mem['h0509] <= 32'hE4E7D8E3;
    mem['h050A] <= 32'h00000013;
    mem['h050B] <= 32'h00000013;
    mem['h050C] <= 32'h02C12083;
    mem['h050D] <= 32'h02812403;
    mem['h050E] <= 32'h03010113;
    mem['h050F] <= 32'h00008067;
    mem['h0510] <= 32'hF4010113;
    mem['h0511] <= 32'h0A112E23;
    mem['h0512] <= 32'h0A812C23;
    mem['h0513] <= 32'h0C010413;
    mem['h0514] <= 32'hF4A42623;
    mem['h0515] <= 32'hF4B42423;
    mem['h0516] <= 32'hF4C42223;
    mem['h0517] <= 32'hF7C40793;
    mem['h0518] <= 32'h00078513;
    mem['h0519] <= 32'h9D9FF0EF;
    mem['h051A] <= 32'hF7C40793;
    mem['h051B] <= 32'hF4842603;
    mem['h051C] <= 32'hF4C42583;
    mem['h051D] <= 32'h00078513;
    mem['h051E] <= 32'hA85FF0EF;
    mem['h051F] <= 32'hF5C40713;
    mem['h0520] <= 32'hF7C40793;
    mem['h0521] <= 32'h00070593;
    mem['h0522] <= 32'h00078513;
    mem['h0523] <= 32'hB81FF0EF;
    mem['h0524] <= 32'hFE042623;
    mem['h0525] <= 32'h0680006F;
    mem['h0526] <= 32'hFEC42783;
    mem['h0527] <= 32'hFF078793;
    mem['h0528] <= 32'h008787B3;
    mem['h0529] <= 32'hF6C7C783;
    mem['h052A] <= 32'hF5840713;
    mem['h052B] <= 32'h00070593;
    mem['h052C] <= 32'h00078513;
    mem['h052D] <= 32'hBC4FF0EF;
    mem['h052E] <= 32'hFEC42783;
    mem['h052F] <= 32'h00179793;
    mem['h0530] <= 32'h00078713;
    mem['h0531] <= 32'hF4442783;
    mem['h0532] <= 32'h00E787B3;
    mem['h0533] <= 32'hF5844703;
    mem['h0534] <= 32'h00E78023;
    mem['h0535] <= 32'hFEC42783;
    mem['h0536] <= 32'h00179793;
    mem['h0537] <= 32'h00178793;
    mem['h0538] <= 32'hF4442703;
    mem['h0539] <= 32'h00F707B3;
    mem['h053A] <= 32'hF5944703;
    mem['h053B] <= 32'h00E78023;
    mem['h053C] <= 32'hFEC42783;
    mem['h053D] <= 32'h00178793;
    mem['h053E] <= 32'hFEF42623;
    mem['h053F] <= 32'hFEC42703;
    mem['h0540] <= 32'h01F00793;
    mem['h0541] <= 32'hF8E7DAE3;
    mem['h0542] <= 32'hF4442783;
    mem['h0543] <= 32'h04078793;
    mem['h0544] <= 32'h00078023;
    mem['h0545] <= 32'h00000013;
    mem['h0546] <= 32'h0BC12083;
    mem['h0547] <= 32'h0B812403;
    mem['h0548] <= 32'h0C010113;
    mem['h0549] <= 32'h00008067;
    mem['h054A] <= 32'h746F6F42;
    mem['h054B] <= 32'h20676E69;
    mem['h054C] <= 32'h6F636950;
    mem['h054D] <= 32'h2E636F53;
    mem['h054E] <= 32'h000A2E2E;
    mem['h054F] <= 32'h73657250;
    mem['h0550] <= 32'h4E452073;
    mem['h0551] <= 32'h20524554;
    mem['h0552] <= 32'h63206F74;
    mem['h0553] <= 32'h69746E6F;
    mem['h0554] <= 32'h2E65756E;
    mem['h0555] <= 32'h000A2E2E;
    mem['h0556] <= 32'h0000000A;
    mem['h0557] <= 32'h5F5F2020;
    mem['h0558] <= 32'h20205F5F;
    mem['h0559] <= 32'h2020205F;
    mem['h055A] <= 32'h20202020;
    mem['h055B] <= 32'h5F202020;
    mem['h055C] <= 32'h205F5F5F;
    mem['h055D] <= 32'h20202020;
    mem['h055E] <= 32'h20202020;
    mem['h055F] <= 32'h5F5F5F5F;
    mem['h0560] <= 32'h0000000A;
    mem['h0561] <= 32'h20207C20;
    mem['h0562] <= 32'h285C205F;
    mem['h0563] <= 32'h5F20295F;
    mem['h0564] <= 32'h5F205F5F;
    mem['h0565] <= 32'h202F5F5F;
    mem['h0566] <= 32'h7C5F5F5F;
    mem['h0567] <= 32'h5F5F2020;
    mem['h0568] <= 32'h2F20205F;
    mem['h0569] <= 32'h5F5F5F20;
    mem['h056A] <= 32'h00000A7C;
    mem['h056B] <= 32'h7C207C20;
    mem['h056C] <= 32'h7C20295F;
    mem['h056D] <= 32'h202F7C20;
    mem['h056E] <= 32'h202F5F5F;
    mem['h056F] <= 32'h5F5C205F;
    mem['h0570] <= 32'h5C205F5F;
    mem['h0571] <= 32'h5F202F20;
    mem['h0572] <= 32'h207C5C20;
    mem['h0573] <= 32'h00000A7C;
    mem['h0574] <= 32'h20207C20;
    mem['h0575] <= 32'h7C2F5F5F;
    mem['h0576] <= 32'h28207C20;
    mem['h0577] <= 32'h28207C5F;
    mem['h0578] <= 32'h7C20295F;
    mem['h0579] <= 32'h20295F5F;
    mem['h057A] <= 32'h5F28207C;
    mem['h057B] <= 32'h207C2029;
    mem['h057C] <= 32'h5F5F5F7C;
    mem['h057D] <= 32'h0000000A;
    mem['h057E] <= 32'h7C5F7C20;
    mem['h057F] <= 32'h7C202020;
    mem['h0580] <= 32'h5F5C7C5F;
    mem['h0581] <= 32'h5F5C5F5F;
    mem['h0582] <= 32'h5F2F5F5F;
    mem['h0583] <= 32'h2F5F5F5F;
    mem['h0584] <= 32'h5F5F5C20;
    mem['h0585] <= 32'h5C202F5F;
    mem['h0586] <= 32'h5F5F5F5F;
    mem['h0587] <= 32'h00000A7C;
    mem['h0588] <= 32'h72617453;
    mem['h0589] <= 32'h676E6974;
    mem['h058A] <= 32'h41485320;
    mem['h058B] <= 32'h3635322D;
    mem['h058C] <= 32'h0A2E2E2E;
    mem['h058D] <= 32'h00000000;
    mem['h058E] <= 32'h2D414853;
    mem['h058F] <= 32'h20363532;
    mem['h0590] <= 32'h656E6F44;
    mem['h0591] <= 32'h00000A21;
    mem['h0592] <= 32'h61746144;
    mem['h0593] <= 32'h0000203A;
    mem['h0594] <= 32'h65676944;
    mem['h0595] <= 32'h203A7473;
    mem['h0596] <= 32'h00000000;
    mem['h0597] <= 32'h6C6C6548;
    mem['h0598] <= 32'h57202C6F;
    mem['h0599] <= 32'h646C726F;
    mem['h059A] <= 32'h00000021;
    mem['h059B] <= 32'h33323130;
    mem['h059C] <= 32'h37363534;
    mem['h059D] <= 32'h62613938;
    mem['h059E] <= 32'h66656463;
    mem['h059F] <= 32'h00000000;
    mem['h05A0] <= 32'h30313D3E;
    mem['h05A1] <= 32'h00003030;
    mem['h05A2] <= 32'h33323130;
    mem['h05A3] <= 32'h37363534;
    mem['h05A4] <= 32'h62613938;
    mem['h05A5] <= 32'h66656463;
    mem['h05A6] <= 32'h00000000;
    mem['h05A7] <= 32'h428A2F98;
    mem['h05A8] <= 32'h71374491;
    mem['h05A9] <= 32'hB5C0FBCF;
    mem['h05AA] <= 32'hE9B5DBA5;
    mem['h05AB] <= 32'h3956C25B;
    mem['h05AC] <= 32'h59F111F1;
    mem['h05AD] <= 32'h923F82A4;
    mem['h05AE] <= 32'hAB1C5ED5;
    mem['h05AF] <= 32'hD807AA98;
    mem['h05B0] <= 32'h12835B01;
    mem['h05B1] <= 32'h243185BE;
    mem['h05B2] <= 32'h550C7DC3;
    mem['h05B3] <= 32'h72BE5D74;
    mem['h05B4] <= 32'h80DEB1FE;
    mem['h05B5] <= 32'h9BDC06A7;
    mem['h05B6] <= 32'hC19BF174;
    mem['h05B7] <= 32'hE49B69C1;
    mem['h05B8] <= 32'hEFBE4786;
    mem['h05B9] <= 32'h0FC19DC6;
    mem['h05BA] <= 32'h240CA1CC;
    mem['h05BB] <= 32'h2DE92C6F;
    mem['h05BC] <= 32'h4A7484AA;
    mem['h05BD] <= 32'h5CB0A9DC;
    mem['h05BE] <= 32'h76F988DA;
    mem['h05BF] <= 32'h983E5152;
    mem['h05C0] <= 32'hA831C66D;
    mem['h05C1] <= 32'hB00327C8;
    mem['h05C2] <= 32'hBF597FC7;
    mem['h05C3] <= 32'hC6E00BF3;
    mem['h05C4] <= 32'hD5A79147;
    mem['h05C5] <= 32'h06CA6351;
    mem['h05C6] <= 32'h14292967;
    mem['h05C7] <= 32'h27B70A85;
    mem['h05C8] <= 32'h2E1B2138;
    mem['h05C9] <= 32'h4D2C6DFC;
    mem['h05CA] <= 32'h53380D13;
    mem['h05CB] <= 32'h650A7354;
    mem['h05CC] <= 32'h766A0ABB;
    mem['h05CD] <= 32'h81C2C92E;
    mem['h05CE] <= 32'h92722C85;
    mem['h05CF] <= 32'hA2BFE8A1;
    mem['h05D0] <= 32'hA81A664B;
    mem['h05D1] <= 32'hC24B8B70;
    mem['h05D2] <= 32'hC76C51A3;
    mem['h05D3] <= 32'hD192E819;
    mem['h05D4] <= 32'hD6990624;
    mem['h05D5] <= 32'hF40E3585;
    mem['h05D6] <= 32'h106AA070;
    mem['h05D7] <= 32'h19A4C116;
    mem['h05D8] <= 32'h1E376C08;
    mem['h05D9] <= 32'h2748774C;
    mem['h05DA] <= 32'h34B0BCB5;
    mem['h05DB] <= 32'h391C0CB3;
    mem['h05DC] <= 32'h4ED8AA4A;
    mem['h05DD] <= 32'h5B9CCA4F;
    mem['h05DE] <= 32'h682E6FF3;
    mem['h05DF] <= 32'h748F82EE;
    mem['h05E0] <= 32'h78A5636F;
    mem['h05E1] <= 32'h84C87814;
    mem['h05E2] <= 32'h8CC70208;
    mem['h05E3] <= 32'h90BEFFFA;
    mem['h05E4] <= 32'hA4506CEB;
    mem['h05E5] <= 32'hBEF9A3F7;
    mem['h05E6] <= 32'hC67178F2;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule
